module uart (
    input   wire                    i_clk
);
    
endmodule: uart