`define FIFO_MODE_SYNC